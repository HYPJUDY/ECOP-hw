`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   10:34:44 06/04/2016
// Design Name:   CACHE
// Module Name:   D:/Computer Organization/Cache/v0/test.v
// Project Name:  v0
// Target Device:  
// Tool versions:  
// Description: 
// ��ʵ��Ҫ��ʵ��Cache������Cache�������ַ�任�߼���Ҳ��Cache����������
// ����ֱ��������ַ�任��CPU��Cache�����ݣ����������������뿼���ȴ������ж�ȡ���ݣ�
// Ȼ���ٽ�����д��Cache�У�֮�󣬽���������CPU����Σ�CPU��Ҫ��洢��д���ݡ�
// Verilog Test Fixture created by ISE for module: CACHE
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test;

	// Inputs
	reg clk; // ϵͳʱ�ӣ����ڼ������������ƵȲ�����
	reg clr; // ϵͳ�������źţ�������洢������������
	reg [31:0] AB; // CPU�����ڴ�ĵ�ַ����ַ���ߣ�
	reg [31:0] DB; // 32λ����ΪDB31..DB0���������ߣ�

	reg MWr; // MWr��Ϊ1��д��Ϊ�����д�ź�
	reg RD; // RD��Ϊ0������ΪCache�Ķ��ź�
	wire hit; // �Ƿ����б�־
	wire [31:0] MD; // ������Cache������
	wire [31:0] D; // Cache��CPU����
	wire MRd; // MRd��Ϊ0������Ϊ����Ķ��ź�
	wire WCT; // дCache����洢���ź�

	// Instantiate the Unit Under Test (UUT)
	CACHE CACHE (
		.AB(AB), 
		.DB(DB), 
		.MWr(MWr), 
		.RD(RD), 
		.hit(hit),
		.clk(clk),
		.clr(clr), 
		.MD(MD), 
		.D(D), 
		.MRd(MRd), 
		.WCT(WCT)
	);
	RAM RAM (
	   .AB(AB),
		.DB(DB),
		.MWr(MWr),
		.MRd(MRd),
		.clk(clk),
		.clr(clr),
		.MD(MD)
	);
	TABLE TABLE (
		.AB(AB),
		.DB(DB),
		.clr(clr),
		.WCT(WCT),
		.MWr(MWr),
		.hit(hit)
	);

	// ��һ����Cache�������
	// 1��Cache ���иõ�ַ���ݣ�ֱ�Ӷ�Cache ��������CPU��
	// 2��Cache ���޸õ�ַ���ݣ������Ӵ洢����ȡ�õ�ַ����д��Cache��Ȼ����CPU��

	// �������޸�Cache�ʹ洢��
	// ���Cache���иõ�ַ�����ݣ����޸ģ�û�о�û�еĸ��ˣ���ͬʱ�޸Ĵ洢���õ�ַ��Ԫ���ݡ�


	initial begin
		// Initialize Inputs
      clk = 0;
		clr = 1;
		// Add stimulus here
		#10;
		clr = 0;
		#10;

		// д����10��ʮ���ƣ�ռ�ĸ��ֽڣ��ĸ���Ԫ���� 
		// CacheΪ�գ�û�иõ�ַ�����ݣ�ֻ�޸Ĵ洢���õ�ַ��Ԫ����
		// �洢���д�0x1��ʼ��ţ�ռ4����Ԫ
		AB = 32'b00000000000000000000000000000001;  
		DB = 10;
		RD = 1;
		MWr = 1;
		#50;

		// д����20�� CacheΪ�գ�û�иõ�ַ�����ݣ�ֻ�޸Ĵ洢���õ�ַ��Ԫ����
		AB = 32'b00000000000000000000000000010010;
		DB = 20;
		RD  = 1;
		MWr = 1;
		#50;

		// д����30�� CacheΪ�գ�û�иõ�ַ�����ݣ�ֻ�޸Ĵ洢���õ�ַ��Ԫ����
		AB = 32'b00000000000001000000000000110000;  // 0x40030
		DB = 30;
		RD = 1;
		MWr = 1;
		#50;

	   // �����ݣ�CacheΪ�գ��޸õ�ַ���ݣ������Ӵ洢����ȡ�õ�ַ����д��Cache��Ȼ����CPU
	   // AB = 32'b00000000000001��14λ�����ţ������λ��һλ��Чλ1����ʮ��λ��������11���浽����洢���ĸ��ݿ���ҵ��ĵ�ַ��Ԫ��
		// 00000000000011��14λ��ţ�0000��4λ�����ڵ�ַ���Ӵ洢����ȡ����30д��cache�ĵ�3��ĵ�0-3����Ԫ����110000��ַ��
		AB = 32'b00000000000001000000000000110000;
		RD = 0;
		MWr = 0;
		#50;

		// �����ݣ�CacheΪ�գ��޸õ�ַ���ݣ������Ӵ洢����ȡ�õ�ַ����д��Cache��Ȼ����CPU
	   // AB = 32'b00000000000000��14λ�����ţ������λ��һλ��Чλ1����ʮ��λ��������1���浽����洢���ĸ��ݿ���ҵ��ĵ�ַ��Ԫ��
		// 00000000000001��14λ��ţ�0010��4λ�����ڵ�ַ���Ӵ洢����ȡ����20д��cache�ĵ�1��ĵ�2-5����Ԫ����10010��ַ��
		AB = 32'b00000000000000000000000000010010;
		RD  = 0;
		MWr = 0;
		#50;

		// д����40�� Cache���иõ�ַ�����ݣ��޸�cache��ͬʱ�޸Ĵ洢���õ�ַ��Ԫ���ݡ�
		AB = 32'b00000000000001000000000000110000;
		DB = 40;
		RD = 1;
		MWr = 1;
		#50;

		// д����50�� Cache��û�иõ�ַ�����ݣ�û�����У�ֻ�޸Ĵ洢���õ�ַ��Ԫ����
		// ���11��ǰ����ͬ������ʱCache��block3�Ѿ����ٶ�Ӧ��ַ0x000c0034������block����������洢����Ҫ��block3����Ӧ�ı�־λ��Ϊ0
		AB = 32'b00000000000011000000000000110100;
		DB = 50;
		MWr = 1;
		RD = 1;
		#50;

		// �����ݣ�Cache ���޸õ�ַ���ݣ������Ӵ洢����ȡ�õ�ַ����д��Cache��Ȼ����CPU��
		AB = 32'b00000000000011000000000000110100;  //read
		MWr = 0;
		RD = 0;
		#50;

		// �����ݣ�Cache ���иõ�ַ���ݣ�ֱ�Ӷ�Cache ��������CPU��
		AB = 32'b00000000000000000000000000010010;  //read
		RD = 0;
		MWr = 0;
		#50;
		
		#50;
	end
   always #5 clk=~clk;
endmodule

